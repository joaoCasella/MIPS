library IEEE;
use IEEE.STD_LOGIC_1164.all; use IEEE.NUMERIC_STD_UNSIGNED.all;

entity testbench is
end;

architecture test of testbench is
  component top
  port(clk, reset:           in     STD_LOGIC;
       writedata, aluout:    buffer STD_LOGIC_VECTOR(31 downto 0);
       memwrite:             buffer STD_LOGIC;
       readdata:             STD_LOGIC_VECTOR(31 downto 0);
       srca:                 STD_LOGIC_VECTOR(31 downto 0);
       srcb:                 STD_LOGIC_VECTOR(31 downto 0);
       zero:                 STD_LOGIC;
       pcsrc:                STD_LOGIC
       );
  end component;
  signal writedata, dataadr:    STD_LOGIC_VECTOR(31 downto 0);
  signal clk, reset,  memwrite: STD_LOGIC;
  signal readdata, srca, srcb:  STD_LOGIC_VECTOR(31 downto 0);
  signal zero, pcsrc:           STD_LOGIC;
begin

  -- instantiate device to be tested
  dut: top port map(clk, reset, writedata, dataadr, memwrite, readdata, srca, srcb, zero, pcsrc);

  -- Generate clock with 10 ns period
  process begin
    clk <= '1';
    wait for 5 ns;
    clk <= '0';
    wait for 5 ns;
  end process;

  -- Generate reset for first two clock cycles
  process begin
    reset <= '1';
    wait for 22 ns;
    reset <= '0';
    wait;
  end process;

  -- check that 7 gets written to address 84 at end of program
  process (clk) begin
    if (clk'event and clk = '0' and memwrite = '1') then
      if (to_integer(dataadr) = 84 and to_integer(writedata) = 7) then
        report "NO ERRORS: Simulation succeeded" severity failure;
      elsif (dataadr /= 80) then
        report "Simulation failed" severity failure;
      end if;
    end if;
  end process;
end;
